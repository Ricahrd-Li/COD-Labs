`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 2019/05/08 21:03:57
// Design Name: 
// Module Name: Display
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////

module Display(  
    input [3:0]y,
    output reg[6:0]x
);
    always @ * begin
        case(y[3:0])
            4'b0000: x = 7'b100_0000; //0
            4'b0001: x = 7'b111_1001;//1001_111;
            4'b0010: x = 7'b010_0100;//0010_010;
            4'b0011: x = 7'b011_0000;//0000_110;//
            4'b0100: x = 7'b001_1001;//1001_100;
            4'b0101: x = 7'b001_0010;//0100_100;
            4'b0110: x = 7'b000_0010;//0100_000;
            4'b0111: x = 7'b111_1000;//0001_111;
            4'b1000: x = 7'b000_0000;//0000_000;
            4'b1001: x = 7'b001_0000;//0000_100;
            4'b1010: x= 7'b000_1000; //A 000_1000        
            4'b1011: x= 7'b000_0011; //b 110_0000
            4'b1100: x= 7'b010_0111; //c 111_0010
            4'b1101: x= 7'b010_0001; //d 100_0010
            4'b1110: x= 7'b000_0110;//E  011_0000
            default: x= 7'b000_1110;//F 011_1000
        endcase
      end
      
endmodule
